`include "alu.v"
`include "branch.v"
`include "decoder.v"
`include "memory.v"
`include "regs.v"

`define CLEAN_DATA

module cpu (
    input         i_clk,
    input         i_rst,
    input         i_valid_i,
    input         i_valid_d,
    input  [31:0] i_data_in_i,
    input  [31:0] i_data_in_d,
    output [31:0] o_addr_i,
    output [31:0] o_addr_d,
    output  [3:0] o_we_d,
    output        o_rd_d,
    output [31:0] o_data_out_d);



    /////////////////////////////////////////////////////////////////////////
    // Pipeline Registers
    /////////////////////////////////////////////////////////////////////////

    // Instruction fetch
    reg  [31:0] if_pc;

    // Instruction decode
    reg  [31:0] id_ret;
    reg  [31:0] id_pc;
    reg  [31:0] id_ir;

    // Execute
    reg  [31:0] ex_rsa_d;
    reg  [31:0] ex_rsb_d;
    reg  [31:0] ex_imm;
    reg  [31:0] ex_pc;
    reg  [31:0] ex_ret;
    reg  [ 4:0] ex_opcode;
    reg  [ 2:0] ex_funct3;
    reg         ex_funct7_4;
    reg         ex_alu_pc;
    reg         ex_alu_imm;
    reg         ex_alu_en;
    reg         ex_ma_wr;
    reg         ex_ma_rd;
    reg  [ 1:0] ex_wb_mux;
    reg  [ 4:0] ex_wb_reg;
    reg         ex_wb_en;

    // Memory Access
    reg  [31:0] ma_rsb_d;
    reg  [31:0] ma_alu;
    reg  [31:0] ma_ret;
    reg  [ 2:0] ma_funct3;
    reg         ma_wr;
    reg         ma_rd;
    reg  [ 4:0] ma_wb_reg;
    reg  [ 1:0] ma_wb_mux;
    reg         ma_wb_en;

    // Write Back
    reg  [31:0] wb_wb_d;
    reg  [ 4:0] wb_wb_reg;
    reg         wb_wb_en;



    /////////////////////////////////////////////////////////////////////////
    // Hazard Detection
    /////////////////////////////////////////////////////////////////////////
    wire hz_data;
    reg  hz_branch;
    wire hz_dat_rsa;
    wire hz_dat_rsb;

    assign hz_dat_rsa = hz_rsa && (rsa != 5'b0000) &&
        ((rsa == ex_wb_reg) || (rsa == ma_wb_reg) || (rsa == wb_wb_reg));
    assign hz_dat_rsb = hz_rsb && (rsb != 5'b0000) &&
        ((rsb == ex_wb_reg) || (rsb == ma_wb_reg) || (rsb == wb_wb_reg));

    assign hz_data = hz_dat_rsa || hz_dat_rsb;


    /////////////////////////////////////////////////////////////////////////
    // Clock Enable
    /////////////////////////////////////////////////////////////////////////
    wire clk_ce;

    assign clk_ce = i_valid_i && i_valid_d;



    /////////////////////////////////////////////////////////////////////////
    // Negative Clock
    /////////////////////////////////////////////////////////////////////////
    wire i_clk_n;

    assign i_clk_n = !i_clk;


    /////////////////////////////////////////////////////////////////////////
    // Program Counter
    /////////////////////////////////////////////////////////////////////////
    wire [31:0] pc_next;
    wire [31:0] pc_mux;

    assign pc_next = if_pc + 32'h4;
    assign pc_mux = (branch_en)? alu_out : pc_next;



    /////////////////////////////////////////////////////////////////////////
    // Instruction Fetch Registers
    /////////////////////////////////////////////////////////////////////////

    always @(posedge i_clk) begin
        if (i_rst) begin
            // Clear on reset
            if_pc <= 32'h0;
            hz_branch <= 0;
        end else begin
            // Clear branch hazard if set
            if (hz_branch) begin
                hz_branch <= 0;
            end
            // Update the pc
            if (clk_ce && (!hz_data || branch_en)) begin
                if_pc <= pc_mux;
                // Set hazard if branch taken
                if (branch_en) begin
                    hz_branch <= 1'b1;
                end
            end
        end
    end



    /////////////////////////////////////////////////////////////////////////
    // Instruction Decode Registers
    /////////////////////////////////////////////////////////////////////////

    always @(posedge i_clk) begin
        if (i_rst) begin
            id_ret <= 0;
            id_pc  <= 0;
            id_ir  <= 0;
        end else if (clk_ce && !hz_data) begin
            id_ret <= pc_next;
            id_pc  <= if_pc;
            id_ir  <= i_data_in_i;
        end
        if (branch_en) begin
            id_ir <= 0;
        end
    end



    /////////////////////////////////////////////////////////////////////////
    // Instruction Decoder
    /////////////////////////////////////////////////////////////////////////
    // verilator lint_off unused
    wire [31:0] immediate;
    wire [ 4:0] opcode;
    wire [ 2:0] funct3;
    wire [ 6:0] funct7;
    wire [ 4:0] rsa;
    wire [ 4:0] rsb;
    wire [ 4:0] rd;
    wire        hz_rsa;
    wire        hz_rsb;
    wire        alu_pc;
    wire        alu_imm;
    wire        alu_en;
    wire        d_wr;
    wire        d_rd;
    wire [ 1:0] wb_mux;
    wire        wb_en;
    // verilator lint_on unused

    decoder decoder_i (
        .i_opcode_in (id_ir),
        .o_immediate (immediate),
        .o_opcode    (opcode),
        .o_funct3    (funct3),
        .o_funct7    (funct7),
        .o_rsa       (rsa),
        .o_rsb       (rsb),
        .o_rd        (rd),
        .o_hz_rsa    (hz_rsa),
        .o_hz_rsb    (hz_rsb),
        .o_alu_pc    (alu_pc),
        .o_alu_imm   (alu_imm),
        .o_alu_en    (alu_en),
        .o_ma_wr     (d_wr),
        .o_ma_rd     (d_rd),
        .o_wb_mux    (wb_mux),
        .o_wb_en     (wb_en)
    );



    /////////////////////////////////////////////////////////////////////////
    // Register set
    /////////////////////////////////////////////////////////////////////////
    wire [31:0] rsa_d;
    wire [31:0] rsb_d;

    regs regs_i (
        .i_clk       (i_clk_n),
        .i_we        (wb_wb_en),
        .i_addr_rd_a (rsa),
        .i_addr_rd_b (rsb),
        .i_addr_wr   (wb_wb_reg),
        .i_dat_wr    (wb_wb_d),
        .o_dat_rd_a  (rsa_d),
        .o_dat_rd_b  (rsb_d)
    );



    /////////////////////////////////////////////////////////////////////////
    // Execute Registers
    /////////////////////////////////////////////////////////////////////////

    always @(posedge i_clk) begin
        if (i_rst || hz_branch || hz_data || branch_en) begin
            ex_rsa_d    <= 0;
            ex_rsb_d    <= 0;
            ex_imm      <= 0;
            ex_pc       <= 0;
            ex_ret      <= 0;
            ex_opcode   <= 0;
            ex_funct3   <= 0;
            ex_funct7_4 <= 0;
            ex_alu_pc   <= 0;
            ex_alu_imm  <= 0;
            ex_alu_en   <= 0;
            ex_ma_wr    <= 0;
            ex_ma_rd    <= 0;
            ex_wb_reg   <= 0;
            ex_wb_mux   <= 0;
            ex_wb_en    <= 0;
        end else if (clk_ce) begin
            ex_rsa_d    <= rsa_d;
            ex_rsb_d    <= rsb_d;
            ex_imm      <= immediate;
            ex_pc       <= id_pc;
            ex_ret      <= id_ret;
            ex_opcode   <= opcode;
            ex_funct3   <= funct3;
            ex_funct7_4 <= funct7[4];
            ex_alu_pc   <= alu_pc;
            ex_alu_imm  <= alu_imm;
            ex_alu_en   <= alu_en;
            ex_ma_wr    <= d_wr;
            ex_ma_rd    <= d_rd;
            ex_wb_reg   <= rd;
            ex_wb_mux   <= wb_mux;
            ex_wb_en    <= wb_en;
        end
    end



    /////////////////////////////////////////////////////////////////////////
    // Branch Conditioner
    /////////////////////////////////////////////////////////////////////////
    wire branch_en;

    branch branch_i (
        .i_dat_a  (ex_rsa_d),
        .i_dat_b  (ex_rsb_d),
        .i_funct3 (ex_funct3),
        .i_opcode (ex_opcode),
        .o_branch_en (branch_en)
    );



    /////////////////////////////////////////////////////////////////////////
    // Arythmetic and Logic Unit
    /////////////////////////////////////////////////////////////////////////
    wire [31:0] alu_a_mux;
    wire [31:0] alu_b_mux;
    wire [31:0] alu_out;

    alu alu_i (
        .i_in_a     (alu_a_mux),
        .i_in_b     (alu_b_mux),
        .i_funct3   (ex_funct3),
        .i_funct7_4 (ex_funct7_4),
        .i_alu_en   (ex_alu_en),
        .i_alu_imm  (ex_alu_imm),
        .o_alu_out  (alu_out)
    );

    assign alu_a_mux = (ex_alu_pc)?  ex_pc  : ex_rsa_d;
    assign alu_b_mux = (ex_alu_imm)? ex_imm : ex_rsb_d;



    /////////////////////////////////////////////////////////////////////////
    // Memory Access Registers
    /////////////////////////////////////////////////////////////////////////

    always @(posedge i_clk) begin
        if (i_rst) begin
            ma_rsb_d  <= 0;
            ma_alu    <= 0;
            ma_ret    <= 0;
            ma_funct3 <= 0;
            ma_wr     <= 0;
            ma_rd     <= 0;
            ma_wb_reg <= 0;
            ma_wb_mux <= 0;
            ma_wb_en  <= 0;
        end else if (clk_ce) begin
            ma_rsb_d  <= ex_rsb_d;
            ma_alu    <= alu_out;
            ma_ret    <= ex_ret;
            ma_funct3 <= ex_funct3;
            ma_wr     <= ex_ma_wr;
            ma_rd     <= ex_ma_rd;
            ma_wb_reg <= ex_wb_reg;
            ma_wb_mux <= ex_wb_mux;
            ma_wb_en  <= ex_wb_en;
        end
    end



    /////////////////////////////////////////////////////////////////////////
    // Data Cache
    /////////////////////////////////////////////////////////////////////////
    wire [31:0] ma_rd_dat;
    wire [31:0] ma_wr_dat;
    wire  [3:0] ma_we;
    wire  [3:0] ma_wr_en;
    wire        ma_rd_en;

    memory memory_i (
        .i_data_rd   (i_data_in_d),
        .i_data_wr   (ma_rsb_d),
        .i_shift     (ma_alu[1:0]),
        .i_length    (ma_funct3[1:0]),
        .i_signed_rd (!ma_funct3[2]),
        .o_data_rd   (ma_rd_dat),
        .o_data_wr   (ma_wr_dat),
        .o_we        (ma_we)
    );

    assign ma_wr_en = ma_we & {4{ma_wr && clk_ce}};
    assign ma_rd_en = ma_rd && clk_ce;



    /////////////////////////////////////////////////////////////////////////
    // Write Back Registers
    /////////////////////////////////////////////////////////////////////////
    wire [31:0] wb_dat_mux;

    always @(posedge i_clk) begin
        if (i_rst) begin
            wb_wb_d   <= 0;
            wb_wb_reg <= 0;
            wb_wb_en  <= 0;
        end else if (clk_ce) begin
            wb_wb_d   <= wb_dat_mux;
            wb_wb_reg <= ma_wb_reg;
            wb_wb_en  <= ma_wb_en;
        end
    end

    assign wb_dat_mux = (ma_wb_mux == 2'b10)? ma_ret :
        (ma_wb_mux == 2'b01)? ma_rd_dat : ma_alu;



    /////////////////////////////////////////////////////////////////////////
    // Output assignment
    /////////////////////////////////////////////////////////////////////////
    assign o_addr_i = if_pc;
    assign o_rd_d = ma_rd_en;
    assign o_we_d = ma_wr_en;

`ifdef CLEAN_DATA
    assign o_addr_d     = (ma_rd_en || |ma_wr_en) ? ma_alu : 0;
    assign o_data_out_d = (ma_rd_en || |ma_wr_en) ? ma_wr_dat : 0;
`else
    assign o_addr_d = ma_alu;
    assign o_data_out_d = ma_wr_dat;
`endif


endmodule
