`include "../config.v"

module alu (
  input         i_clk_n,

  input  [31:0] i_in_a,
  input  [31:0] i_in_b,

  input  [ 2:0] i_funct3,
  input  [ 6:0] i_funct7,
  input         i_alu_en,
  input         i_alu_imm,

  output        o_busy,
  output [31:0] o_alu_out
);


  ///////////////////////////////////////////////////////////////////////////
  // Funct7 decoding
  ///////////////////////////////////////////////////////////////////////////
  wire funct7_5 = (i_funct7 == 7'b0100000);

`ifdef MULDIV_EXTENSION
  wire funct7_0 = (i_funct7 == 7'b0000001);
`endif


  ///////////////////////////////////////////////////////////////////////////
  // Adder/subtractor
  ///////////////////////////////////////////////////////////////////////////
  wire op_subtract = i_alu_en && !i_alu_imm && funct7_5;
  wire [31:0] adder_in_b = (op_subtract) ? ~i_in_b : i_in_b;
  wire [31:0] adder_out = i_in_a + adder_in_b + {31'd0, op_subtract};


`ifdef BARREL_SHIFTER

  ///////////////////////////////////////////////////////////////////////////
  // Barrel Shifter
  ///////////////////////////////////////////////////////////////////////////
  // Barrel shifter works in two stages:
  //  Stage 1: value is rotated (not shifted) by given amount of bits
  //  Stage 2: rotated value is masked to form final value

  // Shifter
  wire [31:0] shift_array [0:31];
  wire [31:0] shift_out = shift_array[shift_amount];
  assign shift_array[0] = i_in_a;
  for (genvar i = 0; i < 31; i = i + 1) begin
    assign shift_array[i+1] = { i_in_a[30-i:0], i_in_a[31:31-i] };
  end

  // Mask
  wire [31:0] shift_mask_array [0:31];
  wire [31:0] shift_mask = shift_mask_array[shift_amount];
  for (genvar i = 0; i < 32; i = i + 1) begin
    assign shift_mask_array[i] = (1 << i) - 1;
  end

  // Busy signal
  wire shift_busy = 0;

  // Operation decoder
  wire op_sll = i_alu_en && (i_funct3 == 3'b001);
  wire op_srl = i_alu_en && (i_funct3 == 3'b101) && !funct7_5;
  wire op_sra = i_alu_en && (i_funct3 == 3'b101) &&  funct7_5;
  wire [4:0] shift_amount = (op_sll) ? i_in_b[4:0] : (5'd0 - i_in_b[4:0]);

  // Shift "postprocessing"
  wire [31:0] shift_sll = shift_out & ~shift_mask;
  wire [31:0] shift_srl = shift_out & shift_mask;
  wire [31:0] shift_sra = shift_srl | (~shift_mask & {32{i_in_a[31]}});

  // Final shift mux
  wire [31:0] shift_result = (|shift_amount) ?
    ((op_sra) ? shift_sra : (op_srl) ? shift_srl : shift_sll) : i_in_a;

`else

  ///////////////////////////////////////////////////////////////////////////
  // Bit Shifter
  ///////////////////////////////////////////////////////////////////////////
  reg [31:0] shift_result = 0;
  reg [ 4:0] shift_amount = 0;
  reg        shift_dir_left = 0;

  always @(posedge i_clk_n) begin

    if (op_shift && shift_amount == 0) begin
      shift_amount   <= i_in_b[4:0];
      shift_result   <= i_in_a;
      shift_dir_left <= op_sll;
    end

    if (shift_amount != 0) begin
      shift_result <= (shift_dir_left) ? shift_left : shift_right;
      shift_amount <= shift_amount - 5'h1;
    end

  end

  // Operation decoder
  wire op_sll   = i_alu_en && (i_funct3 == 3'b001);
  wire op_srl   = i_alu_en && (i_funct3 == 3'b101) && !funct7_5;
  wire op_sra   = i_alu_en && (i_funct3 == 3'b101) &&  funct7_5;
  wire op_shift = op_sll || op_srl || op_sra;

  // Shift signals
  wire [31:0] shift_right = {shift_result[31] && op_sra, shift_result[31:1]};
  wire [31:0] shift_left  = {shift_result[30:0], 1'b0};

  // Busy signal
  wire shift_busy = (shift_amount != 0);

`endif


  ///////////////////////////////////////////////////////////////////////////
  // Logic operators
  ///////////////////////////////////////////////////////////////////////////
  wire [31:0] logic_xor = i_in_a ^ i_in_b;
  wire [31:0] logic_or  = i_in_a | i_in_b;
  wire [31:0] logic_and = i_in_a & i_in_b;


  ///////////////////////////////////////////////////////////////////////////
  // Signed/unsigned comparator
  ///////////////////////////////////////////////////////////////////////////
  wire [31:0] comp   = {31'd0, (  $signed(i_in_a) <   $signed(i_in_b))};
  wire [31:0] comp_u = {31'd0, ($unsigned(i_in_a) < $unsigned(i_in_b))};


  ///////////////////////////////////////////////////////////////////////////
  // Final mux
  ///////////////////////////////////////////////////////////////////////////
  wire [31:0] mux_01 = (i_funct3[0] && i_alu_en) ? shift_result : adder_out;
  wire [31:0] mux_23 = (i_funct3[0] && i_alu_en) ? comp_u       : comp;
  wire [31:0] mux_45 = (i_funct3[0] && i_alu_en) ? shift_result : logic_xor;
  wire [31:0] mux_67 = (i_funct3[0] && i_alu_en) ? logic_and    : logic_or;

  wire [31:0] mux_03 = (i_funct3[1] && i_alu_en) ? mux_23 : mux_01;
  wire [31:0] mux_47 = (i_funct3[1] && i_alu_en) ? mux_67 : mux_45;

  wire [31:0] mux_07 = (i_funct3[2] && i_alu_en) ? mux_47 : mux_03;



  ///////////////////////////////////////////////////////////////////////////
  // Multiplier and divider
  ///////////////////////////////////////////////////////////////////////////
`ifdef MULDIV_EXTENSION

  // Inverted input signals
  wire [31:0] in_a_n = (0 - i_in_a[31:0]);
  wire [31:0] in_b_n = (0 - i_in_b[31:0]);

  // Enable signals
  wire md_enable = funct7_0 && i_alu_en && !i_alu_imm;

  // Sign enable signals
  wire md_m_a_signed = (i_funct3 == 3'b001) || (i_funct3 == 3'b010);
  wire md_m_b_signed = (i_funct3 == 3'b001);
  wire md_d_a_signed = (i_funct3 == 3'b100) || (i_funct3 == 3'b110);
  wire md_d_b_signed = (i_funct3 == 3'b100) || (i_funct3 == 3'b110);
  wire md_sign_a = md_m_a_signed || md_d_a_signed;
  wire md_sign_b = md_m_b_signed || md_d_b_signed;

  // Sign signals
  wire [31:0] md_in_a = (i_in_a[31]) ? in_a_n : i_in_a;
  wire [31:0] md_in_b = (i_in_b[31]) ? in_b_n : i_in_b;
  wire md_m_sign = (md_sign_a && i_in_a[31]) ^ (md_sign_b && i_in_b[31]);
  wire md_div_sign = (md_sign_a && i_in_a[31]) ^ (md_sign_b && i_in_b[31]);
  wire md_rem_sign = (md_sign_a && i_in_a[31]);
  wire md_d_sign = (i_funct3[1]) ? md_rem_sign : md_div_sign;

  // Final inputs
  wire [31:0] md_a = (md_sign_a) ? md_in_a : i_in_a;
  wire [31:0] md_b = (md_sign_b) ? md_in_b : i_in_b;

  // Multiplier
`ifdef FAST_MULTIPLIER

  wire [63:0] md_m_mul = md_a * md_b;
  wire        md_m_busy = 0;

`else

  reg  [63:0] md_m_a_reg = 0;
  reg  [31:0] md_m_b_reg = 0;
  reg  [63:0] md_m_mul = 0;

  always @(posedge i_clk_n) begin
    if (md_m_en && ~|md_m_b_reg) begin
      md_m_a_reg <= { 32'd0, md_a };
      md_m_b_reg <= md_b;
      md_m_mul <= 0;
    end else begin
      if (|md_m_b_reg) begin
        if (md_m_b_reg[0]) begin
          md_m_mul <= md_m_mul + md_m_a_reg;
        end
        md_m_a_reg <= { md_m_a_reg[62:0], 1'b0 };
        md_m_b_reg <= { 1'b0, md_m_b_reg[31:1] };
      end
    end
  end

  wire md_m_busy = |md_m_b_reg;
  wire md_m_en = md_enable && !i_funct3[2];

`endif

  // Multiplier "postprocessing"
  wire [63:0] md_m_q = (md_m_sign) ? (0 - md_m_mul) : md_m_mul;
  wire [31:0] md_mul = (|i_funct3[1:0]) ? md_m_q[63:32] : md_m_q[31:0];

  // Divider
  reg [63:0] md_d_a = 0;
  reg [31:0] md_d_b = 0;
  reg [31:0] md_d_q = 0;
  reg [ 5:0] md_d_cnt = 6'b100000;

  always @(posedge i_clk_n) begin
    if (md_d_en) begin
      md_d_a <= { 32'd0, md_a };
      md_d_b <= md_b;
      md_d_q <= 0;
      md_d_cnt <= 0;
    end

    if (!md_d_cnt[5]) begin
      md_d_cnt <= md_d_cnt + 5'd1;
      md_d_q <= { md_d_q[30:0], div_cmp };

      if (div_cmp) begin
        md_d_a <= { md_d_sub[31:0], md_d_a[30:0], 1'b0 };
      end else begin
        md_d_a <= { md_d_a[62:0], 1'b0 };
      end
    end
  end

  wire [31:0] md_d_sub = md_d_a[62:31] - md_d_b;
  wire        div_cmp = (md_d_a[62:31] >= md_d_b);
  wire        md_d_busy = !md_d_cnt[5];
  wire        md_d_en = md_enable &&  i_funct3[2];

  wire [31:0] md_d_div = md_d_q;
  wire [31:0] md_d_rem = md_d_a[63:32];
  wire [31:0] md_d_res = (i_funct3[1]) ? md_d_rem : md_d_div;
  wire [31:0] md_div = (md_d_sign) ? (0 - md_d_res) : md_d_res;

  // Final mux
  wire        md_busy = md_m_busy || md_d_busy;
  wire [31:0] md_result = (i_funct3[2]) ? md_div : md_mul;

`endif


  ///////////////////////////////////////////////////////////////////////////
  // Output assignment
  ///////////////////////////////////////////////////////////////////////////

`ifdef MULDIV_EXTENSION
  assign o_busy = shift_busy || md_busy;
  assign o_alu_out = (md_enable) ? md_result : mux_07;
`else
  assign o_busy = shift_busy;
  assign o_alu_out = mux_07;
`endif


endmodule
